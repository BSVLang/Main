-- Copyright (c) 2014-2019 Bluespec, Inc.  All Rights Reserved.

package DeepThought where

-- ================================================================
-- Interface declaration

interface DeepThought_IFC =
    getAnswer :: ActionValue  (Int 32)

-- ================================================================
-- Module definition

{-# verilog mkDeepThought #-}

mkDeepThought :: Module  DeepThought_IFC
mkDeepThought =
  module
    interface DeepThought_IFC
        getAnswer = return 42

-- ================================================================
