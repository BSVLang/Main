Shifter_iterative.bsv