-- Copyright (c) 2013-2019 Bluespec, Inc. All Rights Reserved.

package Top
where

-- ================================================================
-- Top module for Mergesort example.
-- Instantiates test driver, mergesort, memory, connects them.
-- Dumps a memory region (unsorted).
-- Starts the test driver, waits for completion
-- Dumps the memory region (sorted).

-- ================================================================
-- Bluespec libraries

import Vector
import FIFOF
import GetPut
import ClientServer
import Connectable

-- ----------------
-- Additional libs

-- None

-- ----------------
-- Project imports

import Utils

import Req_Rsp
import Fabric_Defs

import SoC_Map
import Test_Driver
import Memory_Model
import Mergesort

-- ================================================================
-- Top module

{-# verilog mkTop #-}

mkTop :: Module  Empty
mkTop =
  module
    soc_map     :: SoC_Map_IFC     <- mkSoC_Map
    test_driver :: Test_Driver_IFC <- mkTest_Driver
    mem         :: Memory_IFC      <- mkMemory_Model
    mergesort   :: Mergesort_IFC   <- mkMergesort

    -- Connect modules
    mkConnection  test_driver.bus_ifc    mergesort.config_bus_ifc
    mkConnection  mergesort.mem_bus_ifc  mem.bus_ifc

    -- ----------------
    -- Run the test driver

    rg_step :: Reg  (Bit 3) <- mkReg 0

    rules
        -- Initialize memory and mergesort module
        when (rg_step == 0) ==> do
	    $display  "%0d: Top: Initializing memory [%0h..%0h]"
	              cur_cycle
		      soc_map.m_mem0_controller_addr_base
		      soc_map.m_mem0_controller_addr_size
	    mem.init  soc_map.m_mem0_controller_addr_base  soc_map.m_mem0_controller_addr_size
	    mergesort.init  soc_map.m_accel_0_addr_base
	    rg_step := 1

        -- Dump memory (before sorting)
        when (rg_step == 1) ==> do
	    mem.dump_mem_start  (soc_map.m_mem0_controller_addr_base + sort_start_offset)  n_words
	    rg_step := 2

        -- After dump memory region (unsorted), start test driver
        when ((rg_step == 2) && (not mem.dump_mem_busy)) ==> do
            test_driver.start
	    rg_step := 3

        -- After test driver has finished, dump memory (after sorting)
        when ((rg_step == 3) && (not test_driver.busy)) ==> do
	    mem.dump_mem_start  (soc_map.m_mem0_controller_addr_base + sort_start_offset)  n_words
	    rg_step := 4

        -- After dump memory (sorted), stop
        when ((rg_step == 4) && (not mem.dump_mem_busy)) ==> do
            $finish 0

-- ================================================================
