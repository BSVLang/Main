Counter2_Reg.bsv