// Copyright (c) 2018 Bluespec, Inc.  All Rights Reserved

package Project_Params;

// ================================================================
// BSV library imports

// None

// ================================================================
// Project imports

// None

// ================================================================

typedef 32  Addr_Width;
typedef 8   Data_Width;    // Byte-wide

Integer mem_size = 'h_80_0000;    // 8 MB

// ================================================================

endpackage
