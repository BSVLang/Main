MyFIFOF_Reg.bsv