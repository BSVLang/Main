-- Copyright (c) 2013-2019 Bluespec, Inc. All Rights Reserved

package SoC_Fabric
where

-- ================================================================
-- Defines a SoC Fabric that is a specialization of AXI4_Fabric
-- for this particular SoC.

-- ================================================================
-- Project imports

import AXI4_Types
import AXI4_Fabric

import Fabric_Defs       -- for Wd_Addr, Wd_Data, Wd_User
import Fabric_Req_Rsp
import SoC_Map           -- for Num_Initiators, Num_Targets

-- ================================================================
-- Specialization of parameterized AXI4 fabric for this SoC.

type  SoC_Fabric_IFC = AXI4_Fabric_IFC  Num_Initiators
			                Num_Targets
			                Wd_Id
			                Wd_Addr
			                Wd_Data
			                Wd_User

-- Specialization of parameterized AXI4 interfaces for this SoC

type SoC_Fabric_Initiator_IFC = AXI4_Master_IFC  Wd_Id
                                                 Wd_Addr
					         Wd_Data
					         Wd_User

type SoC_Fabric_Target_IFC    = AXI4_Slave_IFC   Wd_Id
                                                 Wd_Addr
					         Wd_Data
					         Wd_User

-- ================================================================
-- The fabric module, specialized

{-# verilog  mkSoC_Fabric #-}

mkSoC_Fabric :: Module  SoC_Fabric_IFC
mkSoC_Fabric =
  module
    soc_map :: SoC_Map_IFC <- mkSoC_Map

    -- Target address decoder.
    -- Identifies whether a given addr is legal and, if so, which target services it.
    let fn_addr_to_target_num :: Fabric_Addr -> (Bool, Target_Num)
        fn_addr_to_target_num    addr =
            -- Mem 0
            if (   (soc_map.m_mem0_controller_addr_base <= addr)
                && (addr < soc_map.m_mem0_controller_addr_lim)) then
                (True, fromInteger mem0_controller_target_num)

            -- UART 0
            else if (   (soc_map.m_uart_0_addr_base <= addr)
                     && (addr < soc_map.m_uart_0_addr_lim)) then
                (True, fromInteger uart_0_target_num)

            -- Accelerator 0
            else if (   (soc_map.m_accel_0_addr_base <= addr)
                     && (addr < soc_map.m_accel_0_addr_lim)) then
                (True, fromInteger accel_0_target_num)

            else
	        (False, _ )

    soc_fabric :: SoC_Fabric_IFC <- mkAXI4_Fabric  fn_addr_to_target_num

    return soc_fabric

-- ================================================================
